module R_at_B_in_Brow_Bcolumn (
    input [9:0] D11,D12,D13,D14,D15,
    input [9:0] D21,D22,D23,D24,D25,
    input [9:0] D31,D32,D33,D34,D35,
    input [9:0] D41,D42,D43,D44,D45,
    input [9:0] D51,D52,D53,D54,D55,

    output [9:0] R 
);

wire [11:0] R_;
//assign R =   +{2'b0,D22[9:2]} + {2'b0,D24[9:2]} + {2'b0,D44[9:2]} + {2'b0,D42[9:2]}
//             +10'd3*{2'b0,D33[9:2]}
//             -10'd3*{4'b0,D13[9:4]}-10'd3*{4'b0,D53[9:4]}-10'd3*{4'b0,D31[9:4]}-10'd3*{4'b0,D35[9:4]};

assign R_ =   +{2'b0,D22[9:2]} + {2'b0,D24[9:2]} + {2'b0,D44[9:2]} + {2'b0,D42[9:2]}
             +{1'b0,D33[9:1]} + {2'b0,D33[9:2]}
             -({3'b0,D13[9:3]} + {4'b0,D13[9:4]} + {3'b0,D53[9:3]} + {4'b0,D53[9:4]} + {3'b0,D31[9:3]} + {4'b0,D31[9:4]} + {3'b0,D35[9:3]} + {4'b0,D35[9:4]});

assign R = (R_[11] == 1)?10'd0:((R_[10]==1)?10'h3FF:R_[9:0]);

endmodule //R_at_B_in_Brow_Bcolumn